�PNG

   IHDR   8       ���    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   ?PLTE�����C��B��A��?��>��=��<��<��<��;��=��;��>��9��:��6��7��:��9��:
(A,   bKGD �H   sIDAT(ϝ�K�@Pb�!0����Y3�)݂6�Uݦ�<3 **�T��q��S��1���b�\Ѡt��RQ������ɝ�"2S�֧̋��@$ϋ^��ӎ�yѶ}m���r?�}Y�^՗    IEND�B`�