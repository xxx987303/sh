�PNG

   IHDR   8       ���    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   �PLTE�����(��*��0��8��:��4������������������7����������)����6��3����������+��"��5��7��"������-��,��/��2��'��%��$��$��-��1��.��1��/��,��.3�O   bKGD �H   �IDAT(�}���0Dс(�����D���?g��P�e���;D�/Z���t�^�~k0G_�{���N�6�Lg��4FQ�E+��e�Z��K7(�P�D��t@]��Hf�(����%G�K5����4ҷC5R�"c����P�4@���U'v��KKT����(;T�RF�x�Z-�P�Ԡ�i���/UUe��(@5�%W!*o�    IEND�B`�