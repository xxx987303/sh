�PNG

   IHDR   8       ���    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   �PLTE�����(��*��0��8��:��4������������������7����������)����6��3����������+��"��5��7��"������-��,��/��2��'��%��$��$��-��1��.��1��/��,��.3�O   bKGD �H   �IDAT(ύ�m� FQ���KŊ�E�1����m�Z��lχ���x>F�7�D��c�y� �R�ȇ�.�Zo�-n�SX��,`I�K�ܸ�0�Sqb���+n�K/%��ݫG��t��Z֪6�p�f�����a����Q�������iB�f]�}N���� 4.���O�֚m�&/V�.$�%�    IEND�B`�